module geriyazma(input [31:0] amb_cikis_i, // Aritmetik Mantık Biriminin çıkış sinyali alındı
                  output [31:0] sonuc_o);   // alınan sinyal yazdırıldı
assign sonuc_o = amb_cikis_i;
endmodule
